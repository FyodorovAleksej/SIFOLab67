lpm_compare1_inst : lpm_compare1 PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		AgB	 => AgB_sig
	);
