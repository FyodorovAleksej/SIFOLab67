lpm_counter1_inst : lpm_counter1 PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
